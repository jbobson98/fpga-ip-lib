module oled_disp (
    input wire clk,
    input wire rst,
    input wire send,
    inout wire i2c_sda,
    inout wire i2c_scl
);






















endmodule